
module SubBytesQuadTestBench();
   initial begin
      $display("\nRUNNING TESTS FOR BYTE ERROR DETECTION");
      
   end
endmodule // SubBytesQuadTestBench
