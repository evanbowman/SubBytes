
module FFMul4(in, out);
   input      [3:0] in;
   output reg [3:0] out;
   
endmodule // FFMul4
